module 32to1mux;

endmodule;